module banner_sys

