module wocky_cp

import os

