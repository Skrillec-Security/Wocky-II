module config